-- Instanciação dos componentes e o mapeamento de portas.\n
<<instance_name>>: <<COMPONENT_NAME>> port map(<<port1>>=><<portX>>, <<port2>>=><<portY>>);
