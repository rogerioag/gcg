-- Declaração dos sinais.\n
signal <<s_sinal_1>>, <<s_sinal_2>>, <<s_sinal_N>>: <<type>> <<length>>;\n
